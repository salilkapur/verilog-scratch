../counter/counter.srcs/sources_1/new/counter_top.sv