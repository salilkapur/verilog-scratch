../counter/counter.srcs/sources_1/new/counter.sv