../counter/counter.srcs/sources_1/new/display.sv